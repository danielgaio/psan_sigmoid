// arquivo contendo a descricao sitetizavel

`timescale 1ns / 1ps

module psoa_sigmoid (
	input 	logic [15:0] x,
	input 	logic clk,
	output 	logic [15:0] f_x
);
	
	always @ (posedge clk) begin

	end // always

endmodule